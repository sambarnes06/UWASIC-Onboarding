module spi_peripheral (
    input wire nCS,
    input wire clk,
    input wire MOSI,
    input wire, MISO
);